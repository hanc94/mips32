`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/03/2021 09:54:42 AM
// Design Name: 
// Module Name: fuentePC_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fuentePC_tb;
reg SaltoCond;
reg zero;

fuentePC UUT();

initial

    begin
    
    
    
    end

endmodule
